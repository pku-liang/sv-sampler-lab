module generated_module(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, var_20, var_21, var_22, var_23, var_24, var_25, var_26, var_27, var_28, var_29, var_30, var_31, var_32, var_33, var_34, var_35, var_36, var_37, var_38, var_39, var_40, var_41, var_42, var_43, var_44, var_45, var_46, var_47, var_48, var_49, x);
    input [4:0] var_0;
    input [4:0] var_1;
    input [6:0] var_2;
    input [6:0] var_3;
    input [4:0] var_4;
    input [4:0] var_5;
    input [5:0] var_6;
    input [5:0] var_7;
    input [6:0] var_8;
    input [7:0] var_9;
    input [7:0] var_10;
    input [3:0] var_11;
    input [3:0] var_12;
    input [3:0] var_13;
    input [6:0] var_14;
    input [7:0] var_15;
    input [3:0] var_16;
    input [5:0] var_17;
    input [4:0] var_18;
    input [7:0] var_19;
    input [7:0] var_20;
    input [3:0] var_21;
    input [6:0] var_22;
    input [6:0] var_23;
    input [7:0] var_24;
    input [6:0] var_25;
    input [5:0] var_26;
    input [6:0] var_27;
    input [7:0] var_28;
    input [3:0] var_29;
    input [3:0] var_30;
    input [7:0] var_31;
    input [7:0] var_32;
    input [6:0] var_33;
    input [3:0] var_34;
    input [4:0] var_35;
    input [3:0] var_36;
    input [4:0] var_37;
    input [3:0] var_38;
    input [6:0] var_39;
    input [3:0] var_40;
    input [7:0] var_41;
    input [7:0] var_42;
    input [6:0] var_43;
    input [3:0] var_44;
    input [3:0] var_45;
    input [7:0] var_46;
    input [6:0] var_47;
    input [7:0] var_48;
    input [7:0] var_49;
    wire constraint_0, constraint_1, constraint_2, constraint_3, constraint_4, constraint_5, constraint_6, constraint_7, constraint_8, constraint_9, constraint_10, constraint_11, constraint_12, constraint_13, constraint_14, constraint_15, constraint_16, constraint_17, constraint_18, constraint_19, constraint_20, constraint_21, constraint_22, constraint_23, constraint_24, constraint_25, constraint_26, constraint_27, constraint_28, constraint_29, constraint_30, constraint_31, constraint_32, constraint_33, constraint_34, constraint_35, constraint_36, constraint_37, constraint_38, constraint_39, constraint_40, constraint_41, constraint_42, constraint_43, constraint_44, constraint_45, constraint_46, constraint_47, constraint_48, constraint_49;
    output wire x;

    assign constraint_0 = |((var_48 * var_0));
    assign constraint_1 = |((~((var_4 | var_40))));
    assign constraint_2 = |((var_11 * var_16));
    assign constraint_3 = |((var_10 - var_49));
    assign constraint_4 = |(((~(var_34)) + 8'h9));
    assign constraint_5 = |((~((!((var_7 - var_49))))));
    assign constraint_6 = |(((var_37 ^ var_1) && var_47));
    assign constraint_7 = |((8'h9 == 0 ? 0 : (8'hf == 0 ? 0 : var_19 / 8'hf) / 8'h9));
    assign constraint_8 = |(((var_31 & var_37) ^ 8'h72));
    assign constraint_9 = |(((!(var_48)) | 1'h1));
    assign constraint_10 = |((7'hd == 0 ? 0 : var_23 / 7'hd));
    assign constraint_11 = |(((var_8 ^ var_38) && var_39));
    assign constraint_12 = |((var_18 >> 5'h3));
    assign constraint_13 = |((var_3 + 8'h39));
    assign constraint_14 = |(((!(var_36)) + 8'h1));
    assign constraint_15 = |(((var_16 + 8'hd) != 8'h9));
    assign constraint_16 = |(((var_25 & var_43) || var_23));
    assign constraint_17 = |(((~(var_33)) * var_43));
    assign constraint_18 = |(((var_6 * 8'hc) || var_2));
    assign constraint_19 = |(((var_9 >> 8'h4) != 8'h9));
    assign constraint_20 = |(((8'hf == 0 ? 0 : var_32 / 8'hf) * 8'h7));
    assign constraint_21 = |((var_27 >> 7'h0));
    assign constraint_22 = |(((~(var_34)) << 4'h1));
    assign constraint_23 = |((var_23 - 8'h74));
    assign constraint_24 = |((!((var_23 - 8'h79) != 0) || (8'h9f != 0)));
    assign constraint_25 = |((var_37 & var_40));
    assign constraint_26 = |(((!(var_20)) ^ 1'h1));
    assign constraint_27 = |(((~(var_48)) | 8'ha6));
    assign constraint_28 = |(((var_24 - 8'hf9) ^ 8'h10));
    assign constraint_29 = |(((~(var_3)) * var_45));
    assign constraint_30 = |(((!(var_48)) + 8'h1));
    assign constraint_31 = |((var_1 << 5'h2));
    assign constraint_32 = |(((var_12 != 8'h7) && var_49));
    assign constraint_33 = |((!((var_25 & 7'h76))));
    assign constraint_34 = |((var_33 != 8'h1b));
    assign constraint_35 = |(((~(var_8)) | 7'h9));
    assign constraint_36 = |((!((~((var_31 - var_23))))));
    assign constraint_37 = |(((~(var_33)) << 7'h5));
    assign constraint_38 = |((!((4'h6 == 0 ? 0 : var_40 / 4'h6))));
    assign constraint_39 = |(((~(var_37)) | var_1));
    assign constraint_40 = |(((var_20 * 8'h1) || var_41));
    assign constraint_41 = |(((!(var_16)) != var_27));
    assign constraint_42 = |(((var_4 >> 5'h2) - var_33));
    assign constraint_43 = |((var_1 ^ var_36));
    assign constraint_44 = |(((var_25 != 8'h44) || var_2));
    assign constraint_45 = |((~((var_2 ^ var_7))));
    assign constraint_46 = |((var_18 & var_4));
    assign constraint_47 = |(((var_11 + 8'hc) != 8'h54));
    assign constraint_48 = |((1'h1 == 0 ? 0 : (!(var_10)) / 1'h1));
    assign constraint_49 = |(((var_46 & var_37) * var_44));
    assign x = constraint_0 & constraint_1 & constraint_2 & constraint_3 & constraint_4 & constraint_5 & constraint_6 & constraint_7 & constraint_8 & constraint_9 & constraint_10 & constraint_11 & constraint_12 & constraint_13 & constraint_14 & constraint_15 & constraint_16 & constraint_17 & constraint_18 & constraint_19 & constraint_20 & constraint_21 & constraint_22 & constraint_23 & constraint_24 & constraint_25 & constraint_26 & constraint_27 & constraint_28 & constraint_29 & constraint_30 & constraint_31 & constraint_32 & constraint_33 & constraint_34 & constraint_35 & constraint_36 & constraint_37 & constraint_38 & constraint_39 & constraint_40 & constraint_41 & constraint_42 & constraint_43 & constraint_44 & constraint_45 & constraint_46 & constraint_47 & constraint_48 & constraint_49;
endmodule
