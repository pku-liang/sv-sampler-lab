module generated_module("var_0", "var_1", "var_2", "var_3", "var_4");
    input [12:0] "var_0";
    input [12:0] "var_1";
    input [13:0] "var_2";
    input [13:0] "var_3";
    input [7:0] "var_4";

    wire constraint_0 = ~((var_3 << 14'h9));
    wire constraint_1 = ((var_2 - 16'h39dd) + 16'he8c3);
    wire constraint_2 = (!(var_1) ^ 1'h1);
    wire constraint_3 = (~(var_4) / 8'h3);
    wire constraint_4 = (!(var_0) >> 1'h0);
    wire constraint_5 = ((var_2 >> 14'h1) ^ var_1);
    wire constraint_6 = (!(var_0) && var_3);
    wire constraint_7 = ~((~(var_4) * var_4));
endmodule
