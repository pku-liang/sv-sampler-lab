module generated_module(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, var_20, var_21, var_22, var_23, var_24, var_25, var_26, var_27, var_28, var_29, var_30, var_31, var_32, var_33, var_34, var_35, var_36, var_37, var_38, var_39, x);
    input [6:0] var_0;
    input [5:0] var_1;
    input [6:0] var_2;
    input [6:0] var_3;
    input [3:0] var_4;
    input [3:0] var_5;
    input [6:0] var_6;
    input [3:0] var_7;
    input [3:0] var_8;
    input [5:0] var_9;
    input [7:0] var_10;
    input [6:0] var_11;
    input [3:0] var_12;
    input [3:0] var_13;
    input [5:0] var_14;
    input [7:0] var_15;
    input [4:0] var_16;
    input [5:0] var_17;
    input [4:0] var_18;
    input [6:0] var_19;
    input [7:0] var_20;
    input [4:0] var_21;
    input [3:0] var_22;
    input [7:0] var_23;
    input [3:0] var_24;
    input [7:0] var_25;
    input [3:0] var_26;
    input [6:0] var_27;
    input [3:0] var_28;
    input [4:0] var_29;
    input [6:0] var_30;
    input [3:0] var_31;
    input [6:0] var_32;
    input [3:0] var_33;
    input [3:0] var_34;
    input [7:0] var_35;
    input [4:0] var_36;
    input [6:0] var_37;
    input [4:0] var_38;
    input [7:0] var_39;
    wire constraint_0, constraint_1, constraint_2, constraint_3, constraint_4, constraint_5, constraint_6, constraint_7, constraint_8, constraint_9, constraint_10, constraint_11, constraint_12, constraint_13, constraint_14, constraint_15, constraint_16, constraint_17, constraint_18, constraint_19, constraint_20, constraint_21, constraint_22, constraint_23, constraint_24, constraint_25, constraint_26, constraint_27, constraint_28, constraint_29, constraint_30, constraint_31, constraint_32, constraint_33, constraint_34, constraint_35, constraint_36, constraint_37, constraint_38, constraint_39;
    output wire x;

    assign constraint_0 = |((!((~(var_14)) != 0) || (6'h24 != 0)));
    assign constraint_1 = |(((~(var_26)) || var_25));
    assign constraint_2 = |((var_39 | var_24));
    assign constraint_3 = |(((!(var_37 != 0) || (var_30 != 0)) || var_0));
    assign constraint_4 = |(((var_25 / 8'ha) + 8'he6));
    assign constraint_5 = |(((!(var_6 != 0) || (7'h72 != 0)) << 1'h0));
    assign constraint_6 = |(((var_36 + 8'h5) * var_14));
    assign constraint_7 = |(((!(var_23)) | 1'h1));
    assign constraint_8 = |((!(var_6 != 0) || (7'h59 != 0)));
    assign constraint_9 = |((var_25 != 8'hf2));
    assign constraint_10 = |((var_13 - var_28));
    assign constraint_11 = |((!(var_20 != 0) || (var_28 != 0)));
    assign constraint_12 = |((~((var_31 - var_13))));
    assign constraint_13 = |((~((var_21 ^ var_34))));
    assign constraint_14 = |((var_0 ^ var_33));
    assign constraint_15 = |((var_32 & 7'h34));
    assign constraint_16 = |(((~(var_24)) & var_31));
    assign constraint_17 = |((var_9 + 8'h1b));
    assign constraint_18 = |(((var_5 + var_19) + 8'h6f));
    assign constraint_19 = |(((~(var_6)) ^ var_18));
    assign constraint_20 = |((~((var_5 != var_10))));
    assign constraint_21 = |(((~(var_6)) || var_15));
    assign constraint_22 = |((var_1 & var_7));
    assign constraint_23 = |(((var_38 + var_39) || var_1));
    assign constraint_24 = |(((var_12 | 4'hb) && var_11));
    assign constraint_25 = |(((!(var_7 != 0) || (var_4 != 0)) * var_10));
    assign constraint_26 = |((var_14 >> 6'h1));
    assign constraint_27 = |((!(var_9 != 0) || (6'h33 != 0)));
    assign constraint_28 = |(((!(var_17)) + var_12));
    assign constraint_29 = |(((~(var_10)) & var_37));
    assign constraint_30 = |(((var_15 != var_29) >> 1'h0));
    assign constraint_31 = |((!((var_37 - 8'hb))));
    assign constraint_32 = |(((~(var_6)) * var_30));
    assign constraint_33 = |((var_10 && var_19));
    assign constraint_34 = |((~((var_30 != var_35))));
    assign constraint_35 = |((var_20 / 8'h1));
    assign constraint_36 = |((~((var_5 / 4'h1))));
    assign constraint_37 = |((var_3 & var_38));
    assign constraint_38 = |(((var_8 << 4'h0) / 4'h2));
    assign constraint_39 = |(((var_31 || var_4) || var_7));
    wire constraint_40, constraint_41, constraint_42, constraint_43;
    assign constraint_40 = |(8'ha);
    assign constraint_41 = |(8'h1);
    assign constraint_42 = |(4'h1);
    assign constraint_43 = |(4'h2);
    assign x = constraint_0 & constraint_1 & constraint_2 & constraint_3 & constraint_4 & constraint_5 & constraint_6 & constraint_7 & constraint_8 & constraint_9 & constraint_10 & constraint_11 & constraint_12 & constraint_13 & constraint_14 & constraint_15 & constraint_16 & constraint_17 & constraint_18 & constraint_19 & constraint_20 & constraint_21 & constraint_22 & constraint_23 & constraint_24 & constraint_25 & constraint_26 & constraint_27 & constraint_28 & constraint_29 & constraint_30 & constraint_31 & constraint_32 & constraint_33 & constraint_34 & constraint_35 & constraint_36 & constraint_37 & constraint_38 & constraint_39 & constraint_40 & constraint_41 & constraint_42 & constraint_43;
endmodule
