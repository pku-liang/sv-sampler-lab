module generated_module(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, var_20, var_21, var_22, var_23, var_24, var_25, var_26, var_27, var_28, var_29, var_30, var_31, var_32, var_33, var_34);
    input [14:0] var_0;
    input [12:0] var_1;
    input [14:0] var_2;
    input [7:0] var_3;
    input [5:0] var_4;
    input [11:0] var_5;
    input [5:0] var_6;
    input [11:0] var_7;
    input [9:0] var_8;
    input [10:0] var_9;
    input [10:0] var_10;
    input [10:0] var_11;
    input [9:0] var_12;
    input [3:0] var_13;
    input [12:0] var_14;
    input [14:0] var_15;
    input [11:0] var_16;
    input [12:0] var_17;
    input [6:0] var_18;
    input [6:0] var_19;
    input [15:0] var_20;
    input [3:0] var_21;
    input [5:0] var_22;
    input [13:0] var_23;
    input [13:0] var_24;
    input [12:0] var_25;
    input [12:0] var_26;
    input [8:0] var_27;
    input [10:0] var_28;
    input [12:0] var_29;
    input [6:0] var_30;
    input [7:0] var_31;
    input [5:0] var_32;
    input [13:0] var_33;
    input [8:0] var_34;

    wire constraint_0 = ~((~(var_13) * var_6));
    wire constraint_1 = (var_10 != 16'h1a2);
    wire constraint_2 = ((var_3 / 8'h5) - var_21);
    wire constraint_3 = (var_31 | 8'h68);
    wire constraint_4 = (~(var_22) | var_21);
    wire constraint_5 = (var_11 ^ var_3);
    wire constraint_6 = (~(var_24) -> var_32);
    wire constraint_7 = (var_9 << 11'h4);
    wire constraint_8 = ((var_32 + var_21) * 8'hf);
    wire constraint_9 = (!(var_22) || var_1);
    wire constraint_10 = (!(var_26) + 16'h1);
    wire constraint_11 = (var_0 -> var_19);
    wire constraint_12 = (var_12 || var_14);
    wire constraint_13 = (~(var_19) * var_6);
    wire constraint_14 = (var_14 - 16'h160);
    wire constraint_15 = (var_24 || var_10);
    wire constraint_16 = ~((!(var_22) * var_13));
    wire constraint_17 = (!(var_14) || var_23);
    wire constraint_18 = ((var_31 != 8'h5d) * var_32);
    wire constraint_19 = (!(var_2) | 1'h1);
    wire constraint_20 = (var_20 << 16'hd);
    wire constraint_21 = ((var_4 ^ var_22) - var_2);
    wire constraint_22 = !(~((var_6 || var_17)));
    wire constraint_23 = ((var_7 || var_17) || var_11);
    wire constraint_24 = (!(var_16) != 16'h1);
    wire constraint_25 = (var_13 - var_31);
    wire constraint_26 = (var_31 || var_3);
    wire constraint_27 = ((var_18 | 7'h2) * var_32);
    wire constraint_28 = (var_6 >> 6'h3);
    wire constraint_29 = ((var_3 * var_6) << 8'h2);
    wire constraint_30 = (var_19 != var_7);
    wire constraint_31 = (!(var_2) - 16'h0);
    wire constraint_32 = (!(var_13) * var_31);
    wire constraint_33 = ((var_33 -> var_6) + var_34);
    wire constraint_34 = !((~(var_1) >> 13'h2));
endmodule
