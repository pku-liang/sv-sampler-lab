module generated_module(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, var_20, var_21, var_22, var_23, var_24, var_25, var_26, var_27, var_28, var_29, var_30, var_31, var_32, var_33, var_34, x);
    input [14:0] var_0;
    input [12:0] var_1;
    input [14:0] var_2;
    input [7:0] var_3;
    input [5:0] var_4;
    input [11:0] var_5;
    input [5:0] var_6;
    input [11:0] var_7;
    input [9:0] var_8;
    input [10:0] var_9;
    input [10:0] var_10;
    input [10:0] var_11;
    input [9:0] var_12;
    input [3:0] var_13;
    input [12:0] var_14;
    input [14:0] var_15;
    input [11:0] var_16;
    input [12:0] var_17;
    input [6:0] var_18;
    input [6:0] var_19;
    input [15:0] var_20;
    input [3:0] var_21;
    input [5:0] var_22;
    input [13:0] var_23;
    input [13:0] var_24;
    input [12:0] var_25;
    input [12:0] var_26;
    input [8:0] var_27;
    input [10:0] var_28;
    input [12:0] var_29;
    input [6:0] var_30;
    input [7:0] var_31;
    input [5:0] var_32;
    input [13:0] var_33;
    input [8:0] var_34;
    wire constraint_0, constraint_1, constraint_2, constraint_3, constraint_4, constraint_5, constraint_6, constraint_7, constraint_8, constraint_9, constraint_10, constraint_11, constraint_12, constraint_13, constraint_14, constraint_15, constraint_16, constraint_17, constraint_18, constraint_19, constraint_20, constraint_21, constraint_22, constraint_23, constraint_24, constraint_25, constraint_26, constraint_27, constraint_28, constraint_29, constraint_30, constraint_31, constraint_32, constraint_33, constraint_34;
    output wire x;

    assign constraint_0 = |((~(((~(var_13)) * var_6))));
    assign constraint_1 = |((var_10 != 16'h1a2));
    assign constraint_2 = |(((var_3 / 8'h5) - var_21));
    assign constraint_3 = |((var_31 | 8'h68));
    assign constraint_4 = |(((~(var_22)) | var_21));
    assign constraint_5 = |((var_11 ^ var_3));
    assign constraint_6 = |((!((~(var_24)) != 0) || (var_32 != 0)));
    assign constraint_7 = |((var_9 << 11'h4));
    assign constraint_8 = |(((var_32 + var_21) * 8'hf));
    assign constraint_9 = |(((!(var_22)) || var_1));
    assign constraint_10 = |(((!(var_26)) + 16'h1));
    assign constraint_11 = |((!(var_0 != 0) || (var_19 != 0)));
    assign constraint_12 = |((var_12 || var_14));
    assign constraint_13 = |(((~(var_19)) * var_6));
    assign constraint_14 = |((var_14 - 16'h160));
    assign constraint_15 = |((var_24 || var_10));
    assign constraint_16 = |((~(((!(var_22)) * var_13))));
    assign constraint_17 = |(((!(var_14)) || var_23));
    assign constraint_18 = |(((var_31 != 8'h5d) * var_32));
    assign constraint_19 = |(((!(var_2)) | 1'h1));
    assign constraint_20 = |((var_20 << 16'hd));
    assign constraint_21 = |(((var_4 ^ var_22) - var_2));
    assign constraint_22 = |((!((~((var_6 || var_17))))));
    assign constraint_23 = |(((var_7 || var_17) || var_11));
    assign constraint_24 = |(((!(var_16)) != 16'h1));
    assign constraint_25 = |((var_13 - var_31));
    assign constraint_26 = |((var_31 || var_3));
    assign constraint_27 = |(((var_18 | 7'h2) * var_32));
    assign constraint_28 = |((var_6 >> 6'h3));
    assign constraint_29 = |(((var_3 * var_6) << 8'h2));
    assign constraint_30 = |((var_19 != var_7));
    assign constraint_31 = |(((!(var_2)) - 16'h0));
    assign constraint_32 = |(((!(var_13)) * var_31));
    assign constraint_33 = |(((!(var_33 != 0) || (var_6 != 0)) + var_34));
    assign constraint_34 = |((!(((~(var_1)) >> 13'h2))));
    wire constraint_35;
    assign constraint_35 = |(8'h5);
    assign x = constraint_0 & constraint_1 & constraint_2 & constraint_3 & constraint_4 & constraint_5 & constraint_6 & constraint_7 & constraint_8 & constraint_9 & constraint_10 & constraint_11 & constraint_12 & constraint_13 & constraint_14 & constraint_15 & constraint_16 & constraint_17 & constraint_18 & constraint_19 & constraint_20 & constraint_21 & constraint_22 & constraint_23 & constraint_24 & constraint_25 & constraint_26 & constraint_27 & constraint_28 & constraint_29 & constraint_30 & constraint_31 & constraint_32 & constraint_33 & constraint_34 & constraint_35;
endmodule
