module generated_module(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, x);
    input [27:0] var_0;
    input [23:0] var_1;
    input [26:0] var_2;
    input [25:0] var_3;
    input [16:0] var_4;
    input [19:0] var_5;
    input [29:0] var_6;
    input [24:0] var_7;
    input [25:0] var_8;
    input [29:0] var_9;
    input [29:0] var_10;
    input [31:0] var_11;
    input [31:0] var_12;
    input [20:0] var_13;
    input [18:0] var_14;
    input [18:0] var_15;
    input [31:0] var_16;
    input [23:0] var_17;
    input [25:0] var_18;
    input [23:0] var_19;
    wire constraint_0, constraint_1, constraint_2, constraint_3, constraint_4, constraint_5, constraint_6, constraint_7, constraint_8, constraint_9, constraint_10, constraint_11, constraint_12, constraint_13, constraint_14, constraint_15, constraint_16, constraint_17, constraint_18, constraint_19;
    output wire x;

    assign constraint_0 = |((!((var_16 && var_14))));
    assign constraint_1 = |(((!(var_18)) || var_11));
    assign constraint_2 = |(((var_19 + var_9) || var_0));
    assign constraint_3 = |(((~(var_19)) + 32'h1c5d02));
    assign constraint_4 = |(((var_7 != 32'h2fa4c8) + var_10));
    assign constraint_5 = |(((var_18 || var_15) + var_17));
    assign constraint_6 = |((!((~((var_2 && var_14))))));
    assign constraint_7 = |(((var_14 << 19'h7) + var_10));
    assign constraint_8 = |(((var_3 + 32'hcae052) || var_0));
    assign constraint_9 = |((var_11 << 32'h1));
    assign constraint_10 = |((~((!((var_12 | 32'h40f249f3))))));
    assign constraint_11 = |((var_17 != 32'h6f6235));
    assign constraint_12 = |((!((var_7 ^ 25'hd2672d))));
    assign constraint_13 = |((~((var_10 != var_11))));
    assign constraint_14 = |((var_1 | var_17));
    assign constraint_15 = |((!((var_5 - 32'h411a2))));
    assign constraint_16 = |(((!(var_12)) - var_2));
    assign constraint_17 = |((var_4 - 32'h9916));
    assign constraint_18 = |((!(((!(var_6)) != var_19))));
    assign constraint_19 = |((var_1 - var_6));
    assign x = constraint_0 & constraint_1 & constraint_2 & constraint_3 & constraint_4 & constraint_5 & constraint_6 & constraint_7 & constraint_8 & constraint_9 & constraint_10 & constraint_11 & constraint_12 & constraint_13 & constraint_14 & constraint_15 & constraint_16 & constraint_17 & constraint_18 & constraint_19;
endmodule
