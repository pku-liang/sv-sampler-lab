module generated_module(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, x);
    input [15:0] var_0;
    input [21:0] var_1;
    input [3:0] var_2;
    input [27:0] var_3;
    input [18:0] var_4;
    input [17:0] var_5;
    input [18:0] var_6;
    input [13:0] var_7;
    input [15:0] var_8;
    input [28:0] var_9;
    wire constraint_0, constraint_1, constraint_2, constraint_3, constraint_4, constraint_5, constraint_6, constraint_7, constraint_8, constraint_9;
    output wire x;

    assign constraint_0 = |((~((var_2 << 4'h0))));
    assign constraint_1 = |((var_4 && var_1));
    assign constraint_2 = |(((!(var_7)) != var_1));
    assign constraint_3 = |(((~(var_2)) * var_2));
    assign constraint_4 = |(((!(var_5)) || var_3));
    assign constraint_5 = |((var_2 || var_6));
    assign constraint_6 = |((~((var_0 && var_6))));
    assign constraint_7 = |((var_2 / 4'h4));
    assign constraint_8 = |((var_8 ^ 16'hb816));
    assign constraint_9 = |(((var_7 != 32'h37fd) ^ 1'h1));
    wire constraint_10;
    assign constraint_10 = |(4'h4);
    assign x = constraint_0 & constraint_1 & constraint_2 & constraint_3 & constraint_4 & constraint_5 & constraint_6 & constraint_7 & constraint_8 & constraint_9 & constraint_10;
endmodule
