module generated_module(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, var_20, var_21, var_22, var_23, var_24, var_25, var_26, var_27, var_28, var_29, var_30, var_31, var_32, var_33, var_34, var_35, var_36, var_37, var_38, var_39, x);
    input [6:0] var_0;
    input [5:0] var_1;
    input [6:0] var_2;
    input [6:0] var_3;
    input [3:0] var_4;
    input [3:0] var_5;
    input [6:0] var_6;
    input [3:0] var_7;
    input [3:0] var_8;
    input [5:0] var_9;
    input [7:0] var_10;
    input [6:0] var_11;
    input [3:0] var_12;
    input [3:0] var_13;
    input [5:0] var_14;
    input [7:0] var_15;
    input [4:0] var_16;
    input [5:0] var_17;
    input [4:0] var_18;
    input [6:0] var_19;
    input [7:0] var_20;
    input [4:0] var_21;
    input [3:0] var_22;
    input [7:0] var_23;
    input [3:0] var_24;
    input [7:0] var_25;
    input [3:0] var_26;
    input [6:0] var_27;
    input [3:0] var_28;
    input [4:0] var_29;
    input [6:0] var_30;
    input [3:0] var_31;
    input [6:0] var_32;
    input [3:0] var_33;
    input [3:0] var_34;
    input [7:0] var_35;
    input [4:0] var_36;
    input [6:0] var_37;
    input [4:0] var_38;
    input [7:0] var_39;
    wire constraint_0, constraint_1, constraint_2, constraint_3, constraint_4, constraint_5, constraint_6, constraint_7, constraint_8, constraint_9, constraint_10, constraint_11, constraint_12, constraint_13, constraint_14, constraint_15, constraint_16, constraint_17, constraint_18, constraint_19, constraint_20, constraint_21, constraint_22, constraint_23, constraint_24, constraint_25, constraint_26, constraint_27, constraint_28, constraint_29, constraint_30, constraint_31, constraint_32, constraint_33, constraint_34, constraint_35, constraint_36, constraint_37, constraint_38, constraint_39;
    output wire x;

    assign constraint_0 = |(((var_24 ^ var_13) | var_5));
    assign constraint_1 = |(((var_23 ^ var_5) + 8'h1e));
    assign constraint_2 = |(((var_19 / 7'ha) | 7'h4e));
    assign constraint_3 = |((!((var_16 - 8'h13))));
    assign constraint_4 = |(((var_37 * var_33) * 8'h1));
    assign constraint_5 = |((!((~(var_33)) != 0) || (4'he != 0)));
    assign constraint_6 = |((!((!(var_20 != 0) || (8'h8 != 0)) != 0) || (1'h1 != 0)));
    assign constraint_7 = |((!((var_19 ^ 7'h3a) != 0) || (var_27 != 0)));
    assign constraint_8 = |(((var_0 << 7'h4) ^ 7'h59));
    assign constraint_9 = |(((var_6 & var_14) & var_4));
    assign constraint_10 = |((var_33 >> 4'h2));
    assign constraint_11 = |((var_26 && var_36));
    assign constraint_12 = |((var_27 - 8'h56));
    assign constraint_13 = |((var_20 != 8'h11));
    assign constraint_14 = |((!((!((var_7 + 8'hf))))));
    assign constraint_15 = |((~((var_32 - var_12))));
    assign constraint_16 = |(((!(var_21)) - var_3));
    assign constraint_17 = |((~((var_27 - 8'h4e))));
    assign constraint_18 = |(((var_1 / 6'he) || var_7));
    assign constraint_19 = |((!((var_1 || var_24))));
    assign constraint_20 = |((var_22 ^ var_12));
    assign constraint_21 = |(((!(var_21)) + 8'h1));
    assign constraint_22 = |(((var_6 - 8'h3a) && var_28));
    assign constraint_23 = |(((var_34 + var_12) ^ 4'h5));
    assign constraint_24 = |((var_33 | var_7));
    assign constraint_25 = |((var_17 - var_6));
    assign constraint_26 = |((~((var_22 || var_23))));
    assign constraint_27 = |(((var_21 != var_0) && var_31));
    assign constraint_28 = |(((var_18 | 5'h6) || var_11));
    assign constraint_29 = |((var_27 << 7'h4));
    assign constraint_30 = |((var_12 >> 4'h0));
    assign constraint_31 = |(((var_36 / 5'h9) || var_31));
    assign constraint_32 = |((!((!(var_17 != 0) || (var_34 != 0)))));
    assign constraint_33 = |((var_27 != var_4));
    assign constraint_34 = |((!(((~(var_16)) - var_14))));
    assign constraint_35 = |((!((!((var_4 != var_11))))));
    assign constraint_36 = |((!((var_3 & var_24))));
    assign constraint_37 = |(((~(var_20)) | var_8));
    assign constraint_38 = |(((var_0 - 8'h1f) / 8'h7));
    assign constraint_39 = |(((~(var_21)) & var_5));
    wire constraint_40, constraint_41, constraint_42, constraint_43;
    assign constraint_40 = |(7'ha);
    assign constraint_41 = |(6'he);
    assign constraint_42 = |(5'h9);
    assign constraint_43 = |(8'h7);
    assign x = constraint_0 & constraint_1 & constraint_2 & constraint_3 & constraint_4 & constraint_5 & constraint_6 & constraint_7 & constraint_8 & constraint_9 & constraint_10 & constraint_11 & constraint_12 & constraint_13 & constraint_14 & constraint_15 & constraint_16 & constraint_17 & constraint_18 & constraint_19 & constraint_20 & constraint_21 & constraint_22 & constraint_23 & constraint_24 & constraint_25 & constraint_26 & constraint_27 & constraint_28 & constraint_29 & constraint_30 & constraint_31 & constraint_32 & constraint_33 & constraint_34 & constraint_35 & constraint_36 & constraint_37 & constraint_38 & constraint_39 & constraint_40 & constraint_41 & constraint_42 & constraint_43;
endmodule
