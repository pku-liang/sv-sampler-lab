module generated_module(var_0, var_1, var_2, var_3, var_4, var_5, var_6, var_7, var_8, var_9, var_10, var_11, var_12, var_13, var_14, var_15, var_16, var_17, var_18, var_19, var_20, var_21, var_22, var_23, var_24, var_25, var_26, var_27, var_28, var_29, x);
    input [28:0] var_0;
    input [26:0] var_1;
    input [12:0] var_2;
    input [23:0] var_3;
    input [3:0] var_4;
    input [26:0] var_5;
    input [9:0] var_6;
    input [16:0] var_7;
    input [11:0] var_8;
    input [31:0] var_9;
    input [31:0] var_10;
    input [20:0] var_11;
    input [13:0] var_12;
    input [31:0] var_13;
    input [7:0] var_14;
    input [17:0] var_15;
    input [7:0] var_16;
    input [28:0] var_17;
    input [17:0] var_18;
    input [28:0] var_19;
    input [8:0] var_20;
    input [17:0] var_21;
    input [10:0] var_22;
    input [3:0] var_23;
    input [6:0] var_24;
    input [29:0] var_25;
    input [26:0] var_26;
    input [6:0] var_27;
    input [26:0] var_28;
    input [6:0] var_29;
    wire constraint_0, constraint_1, constraint_2, constraint_3, constraint_4, constraint_5, constraint_6, constraint_7, constraint_8, constraint_9, constraint_10, constraint_11, constraint_12, constraint_13, constraint_14, constraint_15, constraint_16, constraint_17, constraint_18, constraint_19, constraint_20, constraint_21, constraint_22, constraint_23, constraint_24, constraint_25, constraint_26, constraint_27, constraint_28, constraint_29;
    output wire x;

    assign constraint_0 = |(((var_17 + 32'hddeb2bd) | var_9));
    assign constraint_1 = |(((~(var_6)) && var_6));
    assign constraint_2 = |((!(var_19 != 0) || (var_12 != 0)));
    assign constraint_3 = |((var_13 ^ var_20));
    assign constraint_4 = |(((~(var_7)) << 17'h4));
    assign constraint_5 = |((!((~(var_19)) != 0) || (var_19 != 0)));
    assign constraint_6 = |(((~(var_13)) != var_7));
    assign constraint_7 = |((var_20 && var_21));
    assign constraint_8 = |(((var_29 | var_24) - var_11));
    assign constraint_9 = |((var_26 - 32'h624db6d));
    assign constraint_10 = |((!((var_29 + 32'h6a) != 0) || (var_23 != 0)));
    assign constraint_11 = |((var_15 && var_21));
    assign constraint_12 = |(((~(var_14)) * var_4));
    assign constraint_13 = |((var_28 >> 27'h19));
    assign constraint_14 = |((!(var_11 != 0) || (21'h5d4ec != 0)));
    assign constraint_15 = |((var_10 | var_23));
    assign constraint_16 = |((var_27 & var_29));
    assign constraint_17 = |((!(((~(var_12)) & var_16))));
    assign constraint_18 = |((var_24 << 7'h1));
    assign constraint_19 = |(((!(var_20)) + var_11));
    assign constraint_20 = |(((var_25 | var_28) != 32'h1ebe5fcd));
    assign constraint_21 = |(((var_7 || var_16) + var_5));
    assign constraint_22 = |((var_18 & 18'h2579));
    assign constraint_23 = |((var_7 || var_20));
    assign constraint_24 = |(((var_27 != var_2) && var_28));
    assign constraint_25 = |(((var_12 || var_14) & 1'h1));
    assign constraint_26 = |((!(var_20 != 0) || (9'h7f != 0)));
    assign constraint_27 = |((var_10 != var_11));
    assign constraint_28 = |((var_28 - 32'h1369340));
    assign constraint_29 = |(((~(var_27)) * var_29));
    wire constraint_30;
    assign x = constraint_0 & constraint_1 & constraint_2 & constraint_3 & constraint_4 & constraint_5 & constraint_6 & constraint_7 & constraint_8 & constraint_9 & constraint_10 & constraint_11 & constraint_12 & constraint_13 & constraint_14 & constraint_15 & constraint_16 & constraint_17 & constraint_18 & constraint_19 & constraint_20 & constraint_21 & constraint_22 & constraint_23 & constraint_24 & constraint_25 & constraint_26 & constraint_27 & constraint_28 & constraint_29;
endmodule
